netcdf test_file {
  (add badness)
}
