netcdf gathered {
dimensions:
	time = 2 ;
	height = 3 ;
	lat = 4 ;
	lon = 5 ;
	p = 6 ;
	list1 = 4 ;
	list2 = 9 ;
	list3 = 14 ;
variables:
	double time(time) ;
		time:standard_name = "time" ;
		time:units = "days since 2000-1-1" ;
	double height(height) ;
		height:standard_name = "height" ;
		height:units = "metres" ;
		height:positive = "up" ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
	int p(p) ;
		p:long_name = "pseudolevel" ;
	double aux0(list1) ;
		aux0:standard_name = "longitude" ;
		aux0:units = "degrees_east" ;
	double aux1(list3) ;
	double aux2(time, list3, p) ;
	double aux3(p, list3, time) ;
	double aux4(p, time, list3) ;
	double aux5(list3, p, time) ;
	double aux6(list3, time) ;
	double aux7(lat) ;
	double aux8(lon, lat) ;
	double aux9(time, height) ;
	int list1(list1) ;
		list1:compress = "lon" ;
	int list2(list2) ;
		list2:compress = "lat lon" ;
	int list3(list3) ;
		list3:compress = "height lat lon" ;
	double temp1(time, height, lat, list1, p) ;
		temp1:long_name = "temp1" ;
		temp1:units = "K" ;
		temp1:coordinates = "aux0 aux7 aux8 aux9" ;
	double temp2(time, height, list2, p) ;
		temp2:long_name = "temp2" ;
		temp2:units = "K" ;
		temp2:coordinates = "aux7 aux8 aux9" ;
	double temp3(time, list3, p) ;
		temp3:long_name = "temp3" ;
		temp3:units = "K" ;
		temp3:coordinates = "aux0 aux1 aux2 aux3 aux4 aux5 aux6 aux7 aux8 aux9" ;

// global attributes:
		:Conventions = "CF-1.8" ;
data:

 time = 31, 60 ;

 height = 0.5, 1.5, 2.5 ;

 lat = -90, -85, -80, -75 ;

 p = 1, 2, 3, 4, 5, 6 ;

 list1 = 0, 1, 3, 4 ;

 list2 = 0, 1, 5, 6, 13, 14, 17, 18, 19 ;

 list3 = 0, 1, 5, 6, 13, 14, 25, 26, 37, 38, 48, 49, 58, 59 ;
}
