netcdf test_file {
dimensions:
	grid_longitude = 9 ;
	bounds2 = 2 ;
	grid_latitude = 10 ;
	atmosphere_hybrid_height_coordinate = 1 ;
variables:
	double grid_longitude_bounds(grid_longitude, bounds2) ;
	double grid_longitude(grid_longitude) ;
		grid_longitude:standard_name = "grid_longitude" ;
		grid_longitude:units = "degrees" ;
		grid_longitude:bounds = "grid_longitude_bounds" ;
	double grid_latitude(grid_latitude) ;
		grid_latitude:standard_name = "grid_latitude" ;
		grid_latitude:units = "degrees" ;
	double bounds(atmosphere_hybrid_height_coordinate, bounds2) ;
		bounds:formula_terms = "orog: surface_altitude a: bounds_1 b: bounds_2" ;
	double atmosphere_hybrid_height_coordinate(atmosphere_hybrid_height_coordinate) ;
		atmosphere_hybrid_height_coordinate:standard_name = "atmosphere_hybrid_height_coordinate" ;
		atmosphere_hybrid_height_coordinate:bounds = "bounds" ;
		atmosphere_hybrid_height_coordinate:formula_terms = "orog: surface_altitude a: a b: b" ;
	int latitude(grid_latitude, grid_longitude) ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degree_N" ;
	int longitude(grid_longitude, grid_latitude) ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degreesE" ;
	string greek_letters(grid_latitude) ;
		greek_letters:standard_name = "greek_letters" ;
	double bounds_1(atmosphere_hybrid_height_coordinate, bounds2) ;
	double a(atmosphere_hybrid_height_coordinate) ;
		a:units = "m" ;
	double bounds_2(atmosphere_hybrid_height_coordinate, bounds2) ;
	double b(atmosphere_hybrid_height_coordinate) ;
	double surface_altitude(grid_longitude, grid_latitude) ;
		surface_altitude:standard_name = "surface_altitude" ;
		surface_altitude:units = "m" ;
	double cell_measure(grid_longitude, grid_latitude) ;
		cell_measure:units = "km 2" ;
	char rotated_latitude_longitude ;
		rotated_latitude_longitude:grid_mapping_name = "rotated_latitude_longitude" ;
		rotated_latitude_longitude:grid_north_pole_latitude = 38. ;
		rotated_latitude_longitude:grid_north_pole_longitude = 190. ;
	double ancillary0(grid_longitude, grid_latitude) ;
		ancillary0:standard_name = "ancillary0" ;
		ancillary0:units = "m.s-1" ;
	double ancillary1(grid_latitude, grid_longitude) ;
		ancillary1:standard_name = "ancillary1" ;
		ancillary1:units = "m.s-1" ;
	double ancillary2(grid_longitude) ;
		ancillary2:standard_name = "ancillary2" ;
		ancillary2:units = "m.s-1" ;
	double ancillary3(grid_latitude) ;
		ancillary3:standard_name = "ancillary3" ;
		ancillary3:units = "m.s-1" ;
	double eastward_wind(atmosphere_hybrid_height_coordinate, grid_latitude, grid_longitude) ;
		eastward_wind:standard_name = "eastward_wind" ;
		eastward_wind:units = "m s-1" ;
		eastward_wind:flag_values = 1LL, 2LL, 4LL ;
		eastward_wind:flag_meanings = "a bb ccc" ;
		eastward_wind:cell_measures = "area: cell_measure" ;
		eastward_wind:coordinates = "latitude longitude greek_letters" ;
		eastward_wind:grid_mapping = "rotated_latitude_longitude" ;
		eastward_wind:ancillary_variables = "ancillary0 ancillary1 ancillary2 ancillary3" ;
		eastward_wind:cell_methods = "grid_longitude: mean grid_latitude: max" ;

// global attributes:
		:Conventions = "CF-1.8" ;
data:

 grid_longitude_bounds =
  19.5, 20.5,
  20.5, 21.5,
  21.5, 22.5,
  22.5, 23.5,
  23.5, 24.5,
  24.5, 25.5,
  25.5, 26.5,
  26.5, 30,
  30, 36 ;

 grid_longitude = 20, 21, 22, 23, 24, 25, 26, 27, 33 ;

 grid_latitude = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9 ;

 bounds =
  1, 2 ;

 atmosphere_hybrid_height_coordinate = 1.5 ;

 latitude =
  -45, -44, -43, -42, -41, -40, -39, -38, -37,
  -36, -35, -34, -33, -32, -31, -30, -29, -28,
  -27, -26, -25, -24, -23, -22, -21, -20, -19,
  -18, -17, -16, -15, -14, -13, -12, -11, -10,
  -9, -8, -7, -6, -5, -4, -3, -2, -1,
  0, 1, 2, 3, 4, 5, 6, 7, 8,
  9, 10, 11, 12, 13, 14, 15, 16, 17,
  18, 19, 20, 21, 22, 23, 24, 25, 26,
  27, 28, 29, 30, 31, 32, 33, 34, 35,
  36, 37, 38, 39, 40, 41, 42, 43, 44 ;

 longitude =
  60, 61, 62, 63, 64, 65, 66, 67, 68, 69,
  70, 71, 72, 73, 74, 75, 76, 77, 78, 79,
  80, 81, 82, 83, 84, 85, 86, 87, 88, 89,
  90, 91, 92, 93, 94, 95, 96, 97, 98, 99,
  100, 101, 102, 103, 104, 105, 106, 107, 108, 109,
  110, 111, 112, 113, 114, 115, 116, 117, 118, 119,
  120, 121, 122, 123, 124, 125, 126, 127, 128, 129,
  130, 131, 132, 133, 134, 135, 136, 137, 138, 139,
  140, 141, 142, 143, 144, 145, 146, 147, 148, 149 ;

 greek_letters = _, "beta", "gamma", "delta", "epsilon", "zeta", "eta", 
    "theta", "iota", "kappa" ;

 bounds_1 =
  5, 15 ;

 a = 10 ;

 bounds_2 =
  14, 26 ;

 b = 20 ;

 surface_altitude =
  0, 18, 36, 54, 72, 90, 108, 126, 144, 162,
  2, 20, 38, 56, 74, 92, 110, 128, 146, 164,
  4, 22, 40, 58, 76, 94, 112, 130, 148, 166,
  6, 24, 42, 60, 78, 96, 114, 132, 150, 168,
  8, 26, 44, 62, 80, 98, 116, 134, 152, 170,
  10, 28, 46, 64, 82, 100, 118, 136, 154, 172,
  12, 30, 48, 66, 84, 102, 120, 138, 156, 174,
  14, 32, 50, 68, 86, 104, 122, 140, 158, 176,
  16, 34, 52, 70, 88, 106, 124, 142, 160, 178 ;

 cell_measure =
  1, 1235, 2469, 3703, 4937, 6171, 7405, 8639, 9873, 11107,
  12341, 13575, 14809, 16043, 17277, 18511, 19745, 20979, 22213, 23447,
  24681, 25915, 27149, 28383, 29617, 30851, 32085, 33319, 34553, 35787,
  37021, 38255, 39489, 40723, 41957, 43191, 44425, 45659, 46893, 48127,
  49361, 50595, 51829, 53063, 54297, 55531, 56765, 57999, 59233, 60467,
  61701, 62935, 64169, 65403, 66637, 67871, 69105, 70339, 71573, 72807,
  74041, 75275, 76509, 77743, 78977, 80211, 81445, 82679, 83913, 85147,
  86381, 87615, 88849, 90083, 91317, 92551, 93785, 95019, 96253, 97487,
  98721, 99955, 101189, 102423, 103657, 104891, 106125, 107359, 108593, 109827 ;

 rotated_latitude_longitude = "" ;

 ancillary0 =
  0, 0.09, 0.18, 0.27, 0.36, 0.45, 0.54, 0.63, 0.72, 0.81,
  0.01, 0.1, 0.19, 0.28, 0.37, 0.46, 0.55, 0.64, 0.73, 0.82,
  0.02, 0.11, 0.2, 0.29, 0.38, 0.47, 0.56, 0.65, 0.74, 0.83,
  0.03, 0.12, 0.21, 0.3, 0.39, 0.48, 0.57, 0.66, 0.75, 0.84,
  0.04, 0.13, 0.22, 0.31, 0.4, 0.49, 0.58, 0.67, 0.76, 0.85,
  0.05, 0.14, 0.23, 0.32, 0.41, 0.5, 0.59, 0.68, 0.77, 0.86,
  0.06, 0.15, 0.24, 0.33, 0.42, 0.51, 0.6, 0.69, 0.78, 0.87,
  0.07, 0.16, 0.25, 0.34, 0.43, 0.52, 0.61, 0.7, 0.79, 0.88,
  0.08, 0.17, 0.26, 0.35, 0.44, 0.53, 0.62, 0.71, 0.8, 0.89 ;

 ancillary1 =
  0, 0.01, 0.02, 0.03, 0.04, 0.05, 0.06, 0.07, 0.08,
  0.09, 0.1, 0.11, 0.12, 0.13, 0.14, 0.15, 0.16, 0.17,
  0.18, 0.19, 0.2, 0.21, 0.22, 0.23, 0.24, 0.25, 0.26,
  0.27, 0.28, 0.29, 0.3, 0.31, 0.32, 0.33, 0.34, 0.35,
  0.36, 0.37, 0.38, 0.39, 0.4, 0.41, 0.42, 0.43, 0.44,
  0.45, 0.46, 0.47, 0.48, 0.49, 0.5, 0.51, 0.52, 0.53,
  0.54, 0.55, 0.56, 0.57, 0.58, 0.59, 0.6, 0.61, 0.62,
  0.63, 0.64, 0.65, 0.66, 0.67, 0.68, 0.69, 0.7, 0.71,
  0.72, 0.73, 0.74, 0.75, 0.76, 0.77, 0.78, 0.79, 0.8,
  0.81, 0.82, 0.83, 0.84, 0.85, 0.86, 0.87, 0.88, 0.89 ;

 ancillary2 = 0, 0.001, 0.002, 0.003, 0.004, 0.005, 0.006, 0.007, 0.008 ;

 ancillary3 = 0, 0.009, 0.018, 0.027, 0.036, 0.045, 0.054, 0.063, 0.072, 0.081 ;

 eastward_wind =
  0, 1, 2, 3, 4, 5, 6, 7, 8,
  9, 10, 11, 12, 13, 14, 15, 16, 17,
  18, 19, 20, 21, 22, 23, 24, 25, 26,
  27, 28, 29, 30, 31, 32, 33, 34, 35,
  36, 37, 38, 39, 40, 41, 42, 43, 44,
  45, 46, 47, 48, 49, 50, 51, 52, 53,
  54, 55, 56, 57, 58, 59, 60, 61, 62,
  63, 64, 65, 66, 67, 68, 69, 70, 71,
  72, 73, 74, 75, 76, 77, 78, 79, 80,
  81, 82, 83, 84, 85, 86, 87, 88, 89 ;
}
